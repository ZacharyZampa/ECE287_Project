module Subkey_Generator(key, subkey0, subkey1, subkey2,subkey3,subkey4,subkey5,subkey6,subkey7,
			subkey8, subkey9, subkey10, subkey11, subkey12, subkey13, subkey14, subkey15, keyCheck);
			
			input [63:0]key;
			output [47:0]subkey0, subkey1, subkey2,subkey3,subkey4,subkey5,subkey6,subkey7,
			subkey8, subkey9, subkey10, subkey11, subkey12, subkey13, subkey14, subkey15;
			output [63:0]keyCheck;
			
			wire [47:0]subkey0, subkey1, subkey2,subkey3,subkey4,subkey5,subkey6,subkey7,
			subkey8, subkey9, subkey10, subkey11, subkey12, subkey13, subkey14, subkey15;
			
			assign keyCheck = {c0[26], key[41], key[38], key[20], 60'h0};
			
			
			// C (left) and D (right)
			wire [27:0]c0, c1, c2, c3, c4, c5, c6, c7, c8, c9, c10, c11, c12, c13, c14, c15, c16;
			wire [27:0]d0, d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16;
				 
				 
		
			// Define c0 and d0 -----------------------------------------------------------------
			assign c0 =	{ key[56], key[48], key[40], key[32], key[24], key[16], key[8], 
							key[0], key[57], key[49], key[41], key[33], key[25], key[17], 
							key[9], key[1], key[58], key[50], key[42], key[34], key[26], 
							key[18], key[10], key[2], key[59], key[51], key[43], key[35] };

				
			assign d0 =	{ key[62], key[54], key[46], key[38], key[30], key[22], key[14], 
							key[6], key[61], key[53], key[45], key[37], key[29], key[21], 
							key[13], key[5], key[60], key[52], key[44], key[36], key[28], 
							key[20], key[12], key[4], key[27], key[19], key[11], key[3] };

			// End Define c0 and d0 -------------------------------------------------------------
			
			
			
			
			
			// Combined c and d and pc2 permutation ---------------------------------------------
			assign subkey0 = {c1[13], c1[16], c1[10], c1[23], c1[0], c1[4], 
				c1[2], c1[27], c1[14], c1[5], c1[20], c1[9], 
				c1[22], c1[18], c1[11], c1[3], c1[25], c1[7], 
				c1[15], c1[6], c1[26], c1[19], c1[12], c1[1], 
				d1[12], d1[23], d1[2], d1[8], d1[18], d1[26], 
				d1[1], d1[11], d1[22], d1[16], d1[4], d1[19], 
				d1[15], d1[20], d1[10], d1[27], d1[5], d1[24], 
				d1[17], d1[13], d1[21], d1[7], d1[0], d1[3] };

			assign subkey1 = {c2[13], c2[16], c2[10], c2[23], c2[0], c2[4], 
				c2[2], c2[27], c2[14], c2[5], c2[20], c2[9], 
				c2[22], c2[18], c2[11], c2[3], c2[25], c2[7], 
				c2[15], c2[6], c2[26], c2[19], c2[12], c2[1], 
				d2[12], d2[23], d2[2], d2[8], d2[18], d2[26], 
				d2[1], d2[11], d2[22], d2[16], d2[4], d2[19], 
				d2[15], d2[20], d2[10], d2[27], d2[5], d2[24], 
				d2[17], d2[13], d2[21], d2[7], d2[0], d2[3] };

			assign subkey2 = {c3[13], c3[16], c3[10], c3[23], c3[0], c3[4], 
				c3[2], c3[27], c3[14], c3[5], c3[20], c3[9], 
				c3[22], c3[18], c3[11], c3[3], c3[25], c3[7], 
				c3[15], c3[6], c3[26], c3[19], c3[12], c3[1], 
				d3[12], d3[23], d3[2], d3[8], d3[18], d3[26], 
				d3[1], d3[11], d3[22], d3[16], d3[4], d3[19], 
				d3[15], d3[20], d3[10], d3[27], d3[5], d3[24], 
				d3[17], d3[13], d3[21], d3[7], d3[0], d3[3] };

			assign subkey3 = {c4[13], c4[16], c4[10], c4[23], c4[0], c4[4], 
				c4[2], c4[27], c4[14], c4[5], c4[20], c4[9], 
				c4[22], c4[18], c4[11], c4[3], c4[25], c4[7], 
				c4[15], c4[6], c4[26], c4[19], c4[12], c4[1], 
				d4[12], d4[23], d4[2], d4[8], d4[18], d4[26], 
				d4[1], d4[11], d4[22], d4[16], d4[4], d4[19], 
				d4[15], d4[20], d4[10], d4[27], d4[5], d4[24], 
				d4[17], d4[13], d4[21], d4[7], d4[0], d4[3] };

			assign subkey4 = {c5[13], c5[16], c5[10], c5[23], c5[0], c5[4], 
				c5[2], c5[27], c5[14], c5[5], c5[20], c5[9], 
				c5[22], c5[18], c5[11], c5[3], c5[25], c5[7], 
				c5[15], c5[6], c5[26], c5[19], c5[12], c5[1], 
				d5[12], d5[23], d5[2], d5[8], d5[18], d5[26], 
				d5[1], d5[11], d5[22], d5[16], d5[4], d5[19], 
				d5[15], d5[20], d5[10], d5[27], d5[5], d5[24], 
				d5[17], d5[13], d5[21], d5[7], d5[0], d5[3] };

			assign subkey5 = {c6[13], c6[16], c6[10], c6[23], c6[0], c6[4], 
				c6[2], c6[27], c6[14], c6[5], c6[20], c6[9], 
				c6[22], c6[18], c6[11], c6[3], c6[25], c6[7], 
				c6[15], c6[6], c6[26], c6[19], c6[12], c6[1], 
				d6[12], d6[23], d6[2], d6[8], d6[18], d6[26], 
				d6[1], d6[11], d6[22], d6[16], d6[4], d6[19], 
				d6[15], d6[20], d6[10], d6[27], d6[5], d6[24], 
				d6[17], d6[13], d6[21], d6[7], d6[0], d6[3] };

			assign subkey6 = {c7[13], c7[16], c7[10], c7[23], c7[0], c7[4], 
				c7[2], c7[27], c7[14], c7[5], c7[20], c7[9], 
				c7[22], c7[18], c7[11], c7[3], c7[25], c7[7], 
				c7[15], c7[6], c7[26], c7[19], c7[12], c7[1], 
				d7[12], d7[23], d7[2], d7[8], d7[18], d7[26], 
				d7[1], d7[11], d7[22], d7[16], d7[4], d7[19], 
				d7[15], d7[20], d7[10], d7[27], d7[5], d7[24], 
				d7[17], d7[13], d7[21], d7[7], d7[0], d7[3] };

			assign subkey7 = {c8[13], c8[16], c8[10], c8[23], c8[0], c8[4], 
				c8[2], c8[27], c8[14], c8[5], c8[20], c8[9], 
				c8[22], c8[18], c8[11], c8[3], c8[25], c8[7], 
				c8[15], c8[6], c8[26], c8[19], c8[12], c8[1], 
				d8[12], d8[23], d8[2], d8[8], d8[18], d8[26], 
				d8[1], d8[11], d8[22], d8[16], d8[4], d8[19], 
				d8[15], d8[20], d8[10], d8[27], d8[5], d8[24], 
				d8[17], d8[13], d8[21], d8[7], d8[0], d8[3] };

			assign subkey8 = {c9[13], c9[16], c9[10], c9[23], c9[0], c9[4], 
				c9[2], c9[27], c9[14], c9[5], c9[20], c9[9], 
				c9[22], c9[18], c9[11], c9[3], c9[25], c9[7], 
				c9[15], c9[6], c9[26], c9[19], c9[12], c9[1], 
				d9[12], d9[23], d9[2], d9[8], d9[18], d9[26], 
				d9[1], d9[11], d9[22], d9[16], d9[4], d9[19], 
				d9[15], d9[20], d9[10], d9[27], d9[5], d9[24], 
				d9[17], d9[13], d9[21], d9[7], d9[0], d9[3] };

			assign subkey9 = {c10[13], c10[16], c10[10], c10[23], c10[0], c10[4], 
				c10[2], c10[27], c10[14], c10[5], c10[20], c10[9], 
				c10[22], c10[18], c10[11], c10[3], c10[25], c10[7], 
				c10[15], c10[6], c10[26], c10[19], c10[12], c10[1], 
				d10[12], d10[23], d10[2], d10[8], d10[18], d10[26], 
				d10[1], d10[11], d10[22], d10[16], d10[4], d10[19], 
				d10[15], d10[20], d10[10], d10[27], d10[5], d10[24], 
				d10[17], d10[13], d10[21], d10[7], d10[0], d10[3] };

			assign subkey10 = {c11[13], c11[16], c11[10], c11[23], c11[0], c11[4], 
				c11[2], c11[27], c11[14], c11[5], c11[20], c11[9], 
				c11[22], c11[18], c11[11], c11[3], c11[25], c11[7], 
				c11[15], c11[6], c11[26], c11[19], c11[12], c11[1], 
				d11[12], d11[23], d11[2], d11[8], d11[18], d11[26], 
				d11[1], d11[11], d11[22], d11[16], d11[4], d11[19], 
				d11[15], d11[20], d11[10], d11[27], d11[5], d11[24], 
				d11[17], d11[13], d11[21], d11[7], d11[0], d11[3] };

			assign subkey11 = {c12[13], c12[16], c12[10], c12[23], c12[0], c12[4], 
				c12[2], c12[27], c12[14], c12[5], c12[20], c12[9], 
				c12[22], c12[18], c12[11], c12[3], c12[25], c12[7], 
				c12[15], c12[6], c12[26], c12[19], c12[12], c12[1], 
				d12[12], d12[23], d12[2], d12[8], d12[18], d12[26], 
				d12[1], d12[11], d12[22], d12[16], d12[4], d12[19], 
				d12[15], d12[20], d12[10], d12[27], d12[5], d12[24], 
				d12[17], d12[13], d12[21], d12[7], d12[0], d12[3] };

			assign subkey12 = {c13[13], c13[16], c13[10], c13[23], c13[0], c13[4], 
				c13[2], c13[27], c13[14], c13[5], c13[20], c13[9], 
				c13[22], c13[18], c13[11], c13[3], c13[25], c13[7], 
				c13[15], c13[6], c13[26], c13[19], c13[12], c13[1], 
				d13[12], d13[23], d13[2], d13[8], d13[18], d13[26], 
				d13[1], d13[11], d13[22], d13[16], d13[4], d13[19], 
				d13[15], d13[20], d13[10], d13[27], d13[5], d13[24], 
				d13[17], d13[13], d13[21], d13[7], d13[0], d13[3] };

			assign subkey13 = {c14[13], c14[16], c14[10], c14[23], c14[0], c14[4], 
				c14[2], c14[27], c14[14], c14[5], c14[20], c14[9], 
				c14[22], c14[18], c14[11], c14[3], c14[25], c14[7], 
				c14[15], c14[6], c14[26], c14[19], c14[12], c14[1], 
				d14[12], d14[23], d14[2], d14[8], d14[18], d14[26], 
				d14[1], d14[11], d14[22], d14[16], d14[4], d14[19], 
				d14[15], d14[20], d14[10], d14[27], d14[5], d14[24], 
				d14[17], d14[13], d14[21], d14[7], d14[0], d14[3] };

			assign subkey14 = {c15[13], c15[16], c15[10], c15[23], c15[0], c15[4], 
				c15[2], c15[27], c15[14], c15[5], c15[20], c15[9], 
				c15[22], c15[18], c15[11], c15[3], c15[25], c15[7], 
				c15[15], c15[6], c15[26], c15[19], c15[12], c15[1], 
				d15[12], d15[23], d15[2], d15[8], d15[18], d15[26], 
				d15[1], d15[11], d15[22], d15[16], d15[4], d15[19], 
				d15[15], d15[20], d15[10], d15[27], d15[5], d15[24], 
				d15[17], d15[13], d15[21], d15[7], d15[0], d15[3] };

			assign subkey15 = {c16[13], c16[16], c16[10], c16[23], c16[0], c16[4], 
				c16[2], c16[27], c16[14], c16[5], c16[20], c16[9], 
				c16[22], c16[18], c16[11], c16[3], c16[25], c16[7], 
				c16[15], c16[6], c16[26], c16[19], c16[12], c16[1], 
				d16[12], d16[23], d16[2], d16[8], d16[18], d16[26], 
				d16[1], d16[11], d16[22], d16[16], d16[4], d16[19], 
				d16[15], d16[20], d16[10], d16[27], d16[5], d16[24], 
				d16[17], d16[13], d16[21], d16[7], d16[0], d16[3] };
			// End Combined c and d and pc2 permutation -----------------------------------------
			
			
			
			
			// Subkey shifters ------------------------------------------------------------------
			Shifter shifted_c0(c0, 1'b0 , c1); // 0 is shift 1, 1 is shift 2
			Shifter shifted_c1(c1, 1'b0 , c2);
			Shifter shifted_c2(c2, 1'b1 , c3);
			Shifter shifted_c3(c3, 1'b1 , c4);
			Shifter shifted_c4(c4, 1'b1 , c5);
			Shifter shifted_c5(c5, 1'b1 , c6);
			Shifter shifted_c6(c6, 1'b1 , c7);
			Shifter shifted_c7(c7, 1'b1 , c8);
			Shifter shifted_c8(c8, 1'b0 , c9);
			Shifter shifted_c9(c9, 1'b1 , c10);
			Shifter shifted_c10(c10, 1'b1 , c11);
			Shifter shifted_c11(c11, 1'b1 , c12);
			Shifter shifted_c12(c12, 1'b1 , c13);
			Shifter shifted_c13(c13, 1'b1 , c14);
			Shifter shifted_c14(c14, 1'b1 , c15);
			Shifter shifted_c15(c15, 1'b0 , c16);
			
			Shifter shifted_d0(d0, 1'b0 , d1); // 0 is shift 1, 1 is shift 2
			Shifter shifted_d1(d1, 1'b0 , d2);
			Shifter shifted_d2(d2, 1'b1 , d3);
			Shifter shifted_d3(d3, 1'b1 , d4);
			Shifter shifted_d4(d4, 1'b1 , d5);
			Shifter shifted_d5(d5, 1'b1 , d6);
			Shifter shifted_d6(d6, 1'b1 , d7);
			Shifter shifted_d7(d7, 1'b1 , d8);
			Shifter shifted_d8(d8, 1'b0 , d9);
			Shifter shifted_d9(d9, 1'b1 , d10);
			Shifter shifted_d10(d10, 1'b1 , d11);
			Shifter shifted_d11(d11, 1'b1 , d12);
			Shifter shifted_d12(d12, 1'b1 , d13);
			Shifter shifted_d13(d13, 1'b1 , d14);
			Shifter shifted_d14(d14, 1'b1 , d15);
			Shifter shifted_d15(d15, 1'b0 , d16);
			// End Subkey shifters ------------------------------------------------------------------
			
			
endmodule
			
module Shifter(subkeyHalf[27:0], shiftSize, shiftedkey[27:0]);
	input [27:0]subkeyHalf;
	input shiftSize;
	output [27:0]shiftedkey;
	reg [27:0]shiftedkey;
	
	always @ (*)
	begin
		if (shiftSize == 1'b1)
			shiftedkey = {subkeyHalf[25:0], subkeyHalf[27:26]}; // shift 2
		else
			shiftedkey = {subkeyHalf[26:0], subkeyHalf[27]};    // shift 1
	end
	
endmodule

			